

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.897 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.31457 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.62674 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 6.791 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 32.8571 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 0.1748 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.80808 LAYER METAL6 ;
    ANTENNAPARTIALCUTAREA 0.1296 LAYER VIA67 ;
    ANTENNAPARTIALMETALAREA 44.252 LAYER METAL7 ;
    ANTENNAPARTIALMETALSIDEAREA 260.746 LAYER METAL7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL7 ; 
    ANTENNAMAXAREACAR 847.025 LAYER METAL7 ;
    ANTENNAMAXSIDEAREACAR 4985.94 LAYER METAL7 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.187 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.89947 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.163 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5964 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 13.752 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 66.3395 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 13.096 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 63.1842 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 440.913 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2134.58 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.825 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.96825 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.452 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.17652 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2761 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 79.8246 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 394.134 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 0.283 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.36123 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 5.552 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.8975 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 14.08 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 67.9172 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 414.759 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2008.78 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[0]
  PIN SO[3] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 13.096 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 63.1842 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1235 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 270.565 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1315.01 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.0015 LAYER VIA56 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.883 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.8696 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 14.818 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 71.467 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 1.2 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 1.534 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 7.57094 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 393.486 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 1909.55 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 3.08547 LAYER VIA67 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 3.86 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.759 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6984 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 19.304 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 93.237 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1573 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 157.019 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 765.541 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.59972 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 1.815 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.92255 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.478 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.114 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9347 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 24.979 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 120.29 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.231732 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 11.62 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 56.0846 LAYER METAL5 ;
    ANTENNAGATEAREA 1.0049 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 145.157 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 703.793 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.05698 LAYER VIA56 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.187 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.89947 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.527 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3473 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 6.594 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 32.1019 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6214 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 44.6229 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 211.301 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 3.889 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.8985 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 40.2032 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 187.596 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.354 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.5151 LAYER METAL3 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 62.5584 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 296.952 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.02849 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 63.9354 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 305.402 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.37132 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 7.192 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7859 LAYER METAL5 ;
    ANTENNAGATEAREA 0.3159 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 86.7021 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 415.519 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.37132 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.861 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.14141 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.37 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7821 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.144 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.9398 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6136 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.1807 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 157.125 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.16002 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 15.286 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 73.9105 LAYER METAL5 ;
    ANTENNAGATEAREA 1.508 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 42.3173 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 206.137 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.16002 LAYER VIA56 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 1.361 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.73881 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 13.2256 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 62.5607 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.303 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0822 LAYER METAL3 ;
    ANTENNAGATEAREA 0.3211 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 26.6264 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 128.217 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.856245 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.944 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.54304 LAYER METAL4 ;
    ANTENNAGATEAREA 0.3211 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.6806 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 157.937 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.968671 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 14.476 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 70.5916 LAYER METAL5 ;
    ANTENNAGATEAREA 8.68661 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 42.6443 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 208.13 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.56007 LAYER VIA56 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.273 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.31313 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 19.9145 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 97.5457 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA34 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.15921 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.682 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0928 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 32.3742 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 157.477 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.68566 LAYER VIA34 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.187 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.89947 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.213 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4569 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2054 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 22.2742 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 108.46 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.351509 LAYER VIA34 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 3.679 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8884 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 11.432 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.3727 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4108 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 32.0477 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 155.58 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.703018 LAYER VIA34 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 0.861 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.014 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.87734 LAYER METAL3 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.919 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.42279 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 27.364 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 131.813 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 171.378 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 827.293 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.54599 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNADIFFAREA 4.19 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.162 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3992 LAYER METAL3 ;
  END framing_error
END SYS_TOP

END LIBRARY
