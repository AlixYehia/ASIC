
// ************************************************************* //
// Author : Ali Yehia Abdelmonem
// Date   : 2024-10-10
// ************************************************************* //

`timescale 1ns/1ps

module RST_SYNC_tb ();


/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////

parameter	CLK_PERIOD = 10;
parameter	NUM_STAGES_tb = 3;

/////////////////////////////////////////////////////////
//////////////////// DUT Signals ////////////////////////
/////////////////////////////////////////////////////////

reg							CLK_tb;
reg							RST_tb;
wire							SYNC_RST_tb;


////////////////////////////////////////////////////////
////////////////// initial block /////////////////////// 
////////////////////////////////////////////////////////

initial 
 begin
    // system functions
 	$dumpfile ("RST_SYNC.vcd");
 	$dumpvars;

 	initialize ();

 	// apply test
 	check(1'b0);

 	#(2*CLK_PERIOD);
 	$stop;

 end


////////////////////////////////////////////////////////
/////////////////////// TASKS //////////////////////////
////////////////////////////////////////////////////////

/////////////// Signals Initialization //////////////////

task initialize;
 begin
 	CLK_tb = 1'b0;
 	RST_tb = 1'b1;
 end
endtask


////////////////// Operation Check ////////////////////

task check;
 input RST_task;
 begin
 	@(negedge CLK_tb)
 	RST_tb = RST_task;
 	#(CLK_PERIOD/3)
 	RST_tb = 1'b1;  // de-assert RST
 	@(posedge CLK_tb)
 	#(NUM_STAGES_tb*CLK_PERIOD) 
 	if (SYNC_RST_tb == 1'b1)
 	 begin
 	 	$display("RST_SYNC Operation Passed");
 	 end
 	else
 	 begin
 	 	$display("RST_SYNC Operation Failed");
 	 end
 end
endtask


////////////////////////////////////////////////////////
////////////////// Clock Generator  ////////////////////
////////////////////////////////////////////////////////

always #(CLK_PERIOD/2) CLK_tb = ~CLK_tb;


////////////////////////////////////////////////////////
////////////////// DUT Instantiation  //////////////////
////////////////////////////////////////////////////////

RST_SYNC #(.NUM_STAGES(NUM_STAGES_tb)) DUT (
	.CLK(CLK_tb),
	.RST(RST_tb),
	.SYNC_RST(SYNC_RST_tb)
	);



endmodule
